module SSP(
    input PCLK,
    input CLEAR_B,
    input PSEL,
    input PWRITE,
    input [7:0] PWDATA,
    input SSPCLKIN,
    input SSPFSSIN,
    input SSPRXD,
    output [7:0] PRDATA,
    output SSPOE_B,
    output SSPTXD,
    output SSPCLKOUT,
    output SSPFSSOUT,
    output SSPTXINTR,
    output SSPRXINTR
    );
	//wire sspclk1;
	//wire sspclk2;
	wire [7:0] TxDATA;
	wire VALID, SENT;
	//LogicClockGenerate LogicClkGen(
		//.CLK(PCLK),
		//.SSPCLKOUT(sspclk1),
		//);
TxFIFO TxFIFO_tester (.PSEL(PSEL), .PWRITE(PWRITE), .PWDATA(PWDATA), .CLEAR_B(CLEAR_B), .PCLK(PCLK), .SENT(SENT), .TxDATA(TxDATA), .SSPTXINTR(SSPTXINTR), .VALID(VALID));
TxLogic TxLogic_tester (.PCLK(PCLK), .CLEAR_B(CLEAR_B), .VALID(VALID),
	.TxDATA(TxDATA),
	//Outputs;
	.SSPOE_B(SSPOE_B),		//Output enable signal
	.SSPTXD(SSPTXD),			//1-bit serial data output
	.SSPFSSOUT(SSPFSSOUT),		//begin the next cycle
	.SSPCLKOUT(SSPCLKOUT),		//twice slower than PCLK
	.SENT(SENT)    );       //A pulse signal generated by state 7 & 8)		

endmodule