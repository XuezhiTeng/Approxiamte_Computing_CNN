/home/ecelrc/students/xteng/vlsi1/lab3/rtl/apr/Nov28run1/gscl45nm.lef